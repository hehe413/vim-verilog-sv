always@(posedge clk or negedge rst_n)
begin
    if(rst_n==1'b0)begin
        
    end
    else begin
        
    end
end
