always@(*)
begin
     
end
